--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:08:54 04/04/2015
-- Design Name:   
-- Module Name:   C:/Users/Angel/PracticasE6/Tarea2/Memoria_ROM/ROM_TB.vhd
-- Project Name:  Memoria_ROM
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: ROM
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY ROM_TB IS


END ROM_TB;
 
ARCHITECTURE behavior OF ROM_TB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT ROM
    PORT(
         clk : IN  std_logic;
         addres : IN  std_logic_vector(7 downto 0);
         data_out : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk_tb : std_logic := '0';
   signal addres_tb : std_logic_vector(7 downto 0) := (others => '0');

 	--Outputs
   signal data_out_tb : std_logic_vector(7 downto 0);

   -- Clock period definitions
   constant clk_period : time := 5 ns;
	
	--data
	constant Long_Dir :natural := 8; --DIRECCIONAMIENTO DE 8 BITS
	constant Long_Dat :natural := 8;	--CHAR_SYZE

	constant Long_Rom : natural := 2**Long_Dir;  --DIRECCIONAMIENTO PARA MEMORIA DE 256 BYTES
	type address_bus is array ( Long_Rom - 1 downto 0) of std_logic_vector ( Long_Dat - 1 downto 0); 
	
	constant address_index : address_bus := --CONTROL MANUAL DE LAS 256 DIRECCIONES
 (0 => "00000000",   1 => "00000001",   2 => "00000010",   3 => "00000011",
  4 => "00000100",   5 => "00000101",   6 => "00000110",   7 => "00000111",
  8 => "00001000",   9 => "00001001",  10 => "00001010",  11 => "00001011", 
 12 => "00001100",  13 => "00001101",  14 => "00001110",  15 => "00001111", 
 16 => "00010000",  17 => "00010001",  18 => "00010010",  19 => "00010011", 
 20 => "00010100",  21 => "00010101",  22 => "00010110",  23 => "00010111", 
 24 => "00011000",  25 => "00011001",  26 => "00011010",  27 => "00011011",
 28 => "00011100",  29 => "00011101",  30 => "00011110",  31 => "00011111",
 32 => "00100000",  33 => "00100001",  34 => "00100010",  35 => "00100011",
 36 => "00100100",  37 => "00100101",  38 => "00100110",  39 => "00100111", 
 40 => "00101000",  41 => "00101001",  42 => "00101010",  43 => "00101011", 
 44 => "00101100",  45 => "00101101",  46 => "00101110",  47 => "00101111",
 48 => "00110000",  49 => "00110001",  50 => "00110010",  51 => "00110011", 
 52 => "00110100",  53 => "00110101",  54 => "00110110",  55 => "00110111", 
 56 => "00111000",  57 => "00111001",  58 => "00111010",  59 => "00111011", 
 60 => "00111100",  61 => "00111101",  62 => "00111110",  63 => "00111111", 
 64 => "01000000",  65 => "01000001",  66 => "01000010",  67 => "01000011",
 68 => "01000100",  69 => "01000101",  70 => "01000110",  71 => "01000111", 
 72 => "01001000",  73 => "01001001",  74 => "01001010",  75 => "01001011", 
 76 => "01001100",  77 => "01001101",  78 => "01001110",  79 => "01001111", 
 80 => "01010000",  81 => "01010001",  82 => "01010010",  83 => "01010011", 
 84 => "01010100",  85 => "01010101",  86 => "01010110",  87 => "01010111",
 88 => "01011000",  89 => "01011001",  90 => "01011010",  91 => "01011011", 
 92 => "01011100",  93 => "01011101",  94 => "01011110",  95 => "01011111",
 96 => "01100000",  97 => "01100001",  98 => "01100010",  99 => "01100011", 
100 => "01100100", 101 => "01100101", 102 => "01100110", 103 => "01100111", 
104 => "01101000", 105 => "01101001", 106 => "01101010", 107 => "01101011", 
108 => "01101100", 109 => "01101101", 110 => "01101110", 111 => "01101111", 
112 => "01110000", 113 => "01110001", 114 => "01110010", 115 => "01110011", 
116 => "01110100", 117 => "01110101", 118 => "01110110", 119 => "01110111", 
120 => "01111000", 121 => "01111001", 122 => "01111010", 123 => "01111011", 
124 => "01111100", 125 => "01111101", 126 => "01111110", 127 => "01111111",
128 => "10000000", 129 => "10000001", 130 => "10000010", 131 => "10000011", 
132 => "10000100", 133 => "10000101", 134 => "10000110", 135 => "10000111", 
136 => "10001000", 137 => "10001001", 138 => "10001010", 139 => "10001011", 
140 => "10001100", 141 => "10001101", 142 => "10001110", 143 => "10001111", 
144 => "10010000", 145 => "10010001", 146 => "10010010", 147 => "10010011",
148 => "10010100", 149 => "10010101", 150 => "10010110", 151 => "10010111", 
152 => "10011000", 153 => "10011001", 154 => "10011010", 155 => "10011011", 
156 => "10011100", 157 => "10011101", 158 => "10011110", 159 => "10011111", 
160 => "10100000", 161 => "10100001", 162 => "10100010", 163 => "10100011", 
164 => "10100100", 165 => "10100101", 166 => "10100110", 167 => "10100111",
168 => "10101000", 169 => "10101001", 170 => "10101010", 171 => "10101011",
172 => "10101100", 173 => "10101101", 174 => "10101110", 175 => "10101111", 
176 => "10110000", 177 => "10110001", 178 => "10110010", 179 => "10110011",
180 => "10110100", 181 => "10110101", 182 => "10110110", 183 => "10110111",
184 => "10111000", 185 => "10111001", 186 => "10111010", 187 => "10111011",
188 => "10111100", 189 => "10111101", 190 => "10111110", 191 => "10111111",
192 => "11000000", 193 => "11000001", 194 => "11000010", 195 => "11000011",
196 => "11000100", 197 => "11000101", 198 => "11000110", 199 => "11000111",
200 => "11001000", 201 => "11001001", 202 => "11001010", 203 => "11001011",
204 => "11001100", 205 => "11001101", 206 => "11001110", 207 => "11001111",
208 => "11010000", 209 => "11010001", 210 => "11010010", 211 => "11010011",
212 => "11010100", 213 => "11010101", 214 => "11010110", 215 => "11010111",
216 => "11011000", 217 => "11011001", 218 => "11011010", 219 => "11011011",
220 => "11011100", 221 => "11011101", 222 => "11011110", 223 => "11011111",
224 => "11100000", 225 => "11100001", 226 => "11100010", 227 => "11100011",
228 => "11100100", 229 => "11100101", 230 => "11100110", 231 => "11100111",
232 => "11101000", 233 => "11101001", 234 => "11101010", 235 => "11101011",
236 => "11101100", 237 => "11101101", 238 => "11101110", 239 => "11101111",
240 => "11110000", 241 => "11110001", 242 => "11110010", 243 => "11110011",
244 => "11110100", 245 => "11110101", 246 => "11110110", 247 => "11110111",
248 => "11111000", 249 => "11111001", 250 => "11111010", 251 => "11111011",
252 => "11111100", 253 => "11111101", 254 => "11111110", 255 => "11111111",
others => "00000000"  
	 );
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: ROM PORT MAP (
          clk 			=> clk_tb,
          addres 		=> addres_tb,
          data_out 	=> data_out_tb
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk_tb <= '0';
		wait for clk_period/2;
		clk_tb <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
		addres_tb <= "00000000"; 
      wait for 2.5 ns;
		
		for i in 0 to (Long_Rom - 1) loop
					addres_tb <= address_index(i);
					wait for clk_period;
		end loop;
	end process stim_proc;
		

END;
