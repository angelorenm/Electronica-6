----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:50:05 03/18/2015 
-- Design Name: 	MEMORIA ROM DE 8 BITS
-- Module Name:    ROM - Behavioral 
-- Project Name: 
-- Target Devices: 	ZYNQ XC7Z010
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use work.rom_components.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ROM is
generic(	Long_Dir :natural :=   8; --Direccionamiento de 8 bits
			Long_Dat :natural :=   8  --Tama�o del bus de datos.
		  );
port( clk 		:in STD_LOGIC;
		addres 	:in STD_LOGIC_VECTOR(Long_Dir-1 downto 0);
		data_out :out STD_LOGIC_VECTOR(Long_Dat-1 downto 0) 
	  );
end ROM;

architecture Behavioral of ROM is

constant Long_ROM : natural := 2**Long_Dir;	--Tama�o de la Memoria
type Memoria is array (Long_Rom - 1 downto 0) of
					STD_LOGIC_VECTOR(Long_Dat-1 downto 0); --Pila de Memoria de 8 bits con 256 direcciones		
	
constant mem : Memoria := --valores 8 bits correspondientes a una onda senoidal
 (0 => "01111111",   1 => "10000010",   2 => "10000101",   3 => "10001000",
  4 => "10001100",   5 => "10001111",   6 => "10010010",   7 => "10010101",
  8 => "10011000",   9 => "10011011",  10 => "10011110",  11 => "10100001", 
 12 => "10100100",  13 => "10100111",  14 => "10101010",  15 => "10101101", 
 16 => "10110000",  17 => "10110011",  18 => "10110110",  19 => "10111001", 
 20 => "10111011",  21 => "10111110",  22 => "11000001",  23 => "11000011", 
 24 => "11000110",  25 => "11001001",  26 => "11001011",  27 => "11001110",
 28 => "11010000",  29 => "11010011",  30 => "11010101",  31 => "11010111",
 32 => "11011001",  33 => "11011100",  34 => "11011110",  35 => "11100000",
 36 => "11100010",  37 => "11100100",  38 => "11100110",  39 => "11101000", 
 40 => "11101001",  41 => "11101011",  42 => "11101101",  43 => "11101110", 
 44 => "11110000",  45 => "11110001",  46 => "11110010",  47 => "11110100",
 48 => "11110101",  49 => "11110110",  50 => "11110111",  51 => "11111000", 
 52 => "11111001",  53 => "11111010",  54 => "11111011",  55 => "11111100", 
 56 => "11111100",  57 => "11111101",  58 => "11111101",  59 => "11111110", 
 60 => "11111110",  61 => "11111110",  62 => "11111110",  63 => "11111110", 
 64 => "11111110",  65 => "11111110",  66 => "11111110",  67 => "11111110",
 68 => "11111110",  69 => "11111101",  70 => "11111101",  71 => "11111100", 
 72 => "11111100",  73 => "11111011",  74 => "11111010",  75 => "11111010", 
 76 => "11111001",  77 => "11111000",  78 => "11110111",  79 => "11110110", 
 80 => "11110100",  81 => "11110011",  82 => "11110010",  83 => "11110000", 
 84 => "11101111",  85 => "11101101",  86 => "11101100",  87 => "11101010",
 88 => "11101000",  89 => "11100111",  90 => "11100101",  91 => "11100011", 
 92 => "11100001",  93 => "11011111",  94 => "11011101",  95 => "11011011",
 96 => "11011000",  97 => "11010110",  98 => "11010100",  99 => "11010001", 
100 => "11001111", 101 => "11001100", 102 => "11001010", 103 => "11000111", 
104 => "11000101", 105 => "11000010", 106 => "10111111", 107 => "10111101", 
108 => "10111010", 109 => "10110111", 110 => "10110100", 111 => "10110001", 
112 => "10101111", 113 => "10101100", 114 => "10101001", 115 => "10100110", 
116 => "10100011", 117 => "10100000", 118 => "10011101", 119 => "10011010", 
120 => "10010110", 121 => "10010011", 122 => "10010000", 123 => "10001101", 
124 => "10001010", 125 => "10000111", 126 => "10000100", 127 => "10000001",
128 => "01111101", 129 => "01111010", 130 => "01110111", 131 => "01110100", 
132 => "01110001", 133 => "01101110", 134 => "01101011", 135 => "01101000", 
136 => "01100100", 137 => "01100001", 138 => "01011110", 139 => "01011011", 
140 => "01011000", 141 => "01010101", 142 => "01010010", 143 => "01001111", 
144 => "01001101", 145 => "01001010", 146 => "01000111", 147 => "01000100",
148 => "01000001", 149 => "00111111", 150 => "00111100", 151 => "00111001", 
152 => "00110111", 153 => "00110100", 154 => "00110010", 155 => "00101111", 
156 => "00101101", 157 => "00101010", 158 => "00101000", 159 => "00100110", 
160 => "00100011", 161 => "00100001", 162 => "00011111", 163 => "00011101", 
164 => "00011011", 165 => "00011001", 166 => "00010111", 167 => "00010110",
168 => "00010100", 169 => "00010010", 170 => "00010001", 171 => "00001111",
172 => "00001110", 173 => "00001100", 174 => "00001011", 175 => "00001010", 
176 => "00001000", 177 => "00000111", 178 => "00000110", 179 => "00000101",
180 => "00000100", 181 => "00000100", 182 => "00000011", 183 => "00000010",
184 => "00000010", 185 => "00000001", 186 => "00000001", 187 => "00000000",
188 => "00000000", 189 => "00000000", 190 => "00000000", 191 => "00000000",
192 => "00000000", 193 => "00000000", 194 => "00000000", 195 => "00000000",
196 => "00000000", 197 => "00000001", 198 => "00000001", 199 => "00000010",
200 => "00000010", 201 => "00000011", 202 => "00000100", 203 => "00000101",
204 => "00000110", 205 => "00000111", 206 => "00001000", 207 => "00001001",
208 => "00001010", 209 => "00001100", 210 => "00001101", 211 => "00001110",
212 => "00010000", 213 => "00010001", 214 => "00010011", 215 => "00010101",
216 => "00010110", 217 => "00011000", 218 => "00011010", 219 => "00011100",
220 => "00011110", 221 => "00100000", 222 => "00100010", 223 => "00100101",
224 => "00100111", 225 => "00101001", 226 => "00101011", 227 => "00101110",
228 => "00110000", 229 => "00110011", 230 => "00110101", 231 => "00111000",
232 => "00111011", 233 => "00111101", 234 => "01000000", 235 => "01000011",
236 => "01000101", 237 => "01001000", 238 => "01001011", 239 => "01001110",
240 => "01010001", 241 => "01010100", 242 => "01010111", 243 => "01011010",
244 => "01011101", 245 => "01100000", 246 => "01100011", 247 => "01100110",
248 => "01101001", 249 => "01101100", 250 => "01101111", 251 => "01110010",
252 => "01110110", 253 => "01111001", 254 => "01111100", 255 => "01111111",
others => "00000000"  
	 );

 attribute rom_style: string;
 attribute rom_style of data_out: signal is "block";

BEGIN
	ROM_MEM : process(clk)
	BEGIN
			if rising_edge(clk) then
				data_out <= mem(to_integer(unsigned(addres)));
			end if;
	end process ROM_MEM;
	

end architecture Behavioral;

